module NanoProcessor();

endmodule
