module NanoProcessor(
  input clock,
  output [8:0] gpio);

endmodule
